module PE (
  input [31:0] src1,
  input [31:0] src2,
  input [31:0] inst,
  output reg [31:0] out1
);
  //br
  src1 + src2
  fsrc1 + fsrc2
  fsrc1 * fsrc2
  //load
  //store
  //getelementptr
  //icmp
  //phi
  //call
endmodule
